module test_alu



endmodule
